// Created by ihdl
module sineDecoder (
	input	[6:0] A,
	output reg 	[32:0] Y
);

	always @ (A) begin
		case (A)
			7'b0000000: Y = 33'b000000000000000000000000000000001;
			7'b0000001: Y = 33'b000000000000000000000000000000010;
			7'b0000010: Y = 33'b000000000000000000000000000000100;
			7'b0000011: Y = 33'b000000000000000000000000000000101;
			7'b0000100: Y = 33'b000000000000000000000000000000111;
			7'b0000101: Y = 33'b000000000000000000000000000001101;
			7'b0000110: Y = 33'b000000000000000000000000000001110;
			7'b0000111: Y = 33'b000000000000000000000000000011100;
			7'b0001000: Y = 33'b000000000000000000000000000011101;
			7'b0001001: Y = 33'b000000000000000000000000000011111;
			7'b0001010: Y = 33'b000000000000000000000000000111100;
			7'b0001011: Y = 33'b000000000000000000000000000111110;
			7'b0001100: Y = 33'b000000000000000000000000000111111;
			7'b0001101: Y = 33'b000000000000000000000000001111101;
			7'b0001110: Y = 33'b000000000000000000000000001111110;
			7'b0001111: Y = 33'b000000000000000000000000011111100;
			7'b0010000: Y = 33'b000000000000000000000000011111110;
			7'b0010001: Y = 33'b000000000000000000000000011111111;
			7'b0010010: Y = 33'b000000000000000000000000111111101;
			7'b0010011: Y = 33'b000000000000000000000000111111110;
			7'b0010100: Y = 33'b000000000000000000000001111111100;
			7'b0010101: Y = 33'b000000000000000000000001111111101;
			7'b0010110: Y = 33'b000000000000000000000001111111111;
			7'b0010111: Y = 33'b000000000000000000000011111111100;
			7'b0011000: Y = 33'b000000000000000000000011111111110;
			7'b0011001: Y = 33'b000000000000000000000011111111111;
			7'b0011010: Y = 33'b000000000000000000000111111111101;
			7'b0011011: Y = 33'b000000000000000000000111111111110;
			7'b0011100: Y = 33'b000000000000000000001111111111100;
			7'b0011101: Y = 33'b000000000000000000001111111111101;
			7'b0011110: Y = 33'b000000000000000000001111111111110;
			7'b0011111: Y = 33'b000000000000000000011111111111100;
			7'b0100000: Y = 33'b000000000000000000011111111111101;
			7'b0100001: Y = 33'b000000000000000000011111111111111;
			7'b0100010: Y = 33'b000000000000000000111111111111100;
			7'b0100011: Y = 33'b000000000000000000111111111111110;
			7'b0100100: Y = 33'b000000000000000000111111111111111;
			7'b0100101: Y = 33'b000000000000000001111111111111100;
			7'b0100110: Y = 33'b000000000000000001111111111111110;
			7'b0100111: Y = 33'b000000000000000001111111111111111;
			7'b0101000: Y = 33'b000000000000000011111111111111101;
			7'b0101001: Y = 33'b000000000000000011111111111111110;
			7'b0101010: Y = 33'b000000000000000011111111111111111;
			7'b0101011: Y = 33'b000000000000000111111111111111101;
			7'b0101100: Y = 33'b000000000000000111111111111111110;
			7'b0101101: Y = 33'b000000000000000111111111111111111;
			7'b0101110: Y = 33'b000000000000001111111111111111101;
			7'b0101111: Y = 33'b000000000000001111111111111111110;
			7'b0110000: Y = 33'b000000000000001111111111111111111;
			7'b0110001: Y = 33'b000000000000011111111111111111100;
			7'b0110010: Y = 33'b000000000000011111111111111111110;
			7'b0110011: Y = 33'b000000000000011111111111111111111;
			7'b0110100: Y = 33'b000000000000111111111111111111100;
			7'b0110101: Y = 33'b000000000000111111111111111111110;
			7'b0110110: Y = 33'b000000000000111111111111111111111;
			7'b0110111: Y = 33'b000000000001111111111111111111100;
			7'b0111000: Y = 33'b000000000001111111111111111111101;
			7'b0111001: Y = 33'b000000000001111111111111111111110;
			7'b0111010: Y = 33'b000000000011111111111111111111100;
			7'b0111011: Y = 33'b000000000011111111111111111111101;
			7'b0111100: Y = 33'b000000000011111111111111111111110;
			7'b0111101: Y = 33'b000000000011111111111111111111111;
			7'b0111110: Y = 33'b000000000111111111111111111111100;
			7'b0111111: Y = 33'b000000000111111111111111111111101;
			7'b1000000: Y = 33'b000000000111111111111111111111110;
			7'b1000001: Y = 33'b000000000111111111111111111111111;
			7'b1000010: Y = 33'b000000001111111111111111111111101;
			7'b1000011: Y = 33'b000000001111111111111111111111110;
			7'b1000100: Y = 33'b000000001111111111111111111111111;
			7'b1000101: Y = 33'b000000011111111111111111111111100;
			7'b1000110: Y = 33'b000000011111111111111111111111101;
			7'b1000111: Y = 33'b000000011111111111111111111111110;
			7'b1001000: Y = 33'b000000011111111111111111111111111;
			7'b1001001: Y = 33'b000000111111111111111111111111100;
			7'b1001010: Y = 33'b000000111111111111111111111111101;
			7'b1001011: Y = 33'b000000111111111111111111111111110;
			7'b1001100: Y = 33'b000000111111111111111111111111110;
			7'b1001101: Y = 33'b000000111111111111111111111111111;
			7'b1001110: Y = 33'b000001111111111111111111111111100;
			7'b1001111: Y = 33'b000001111111111111111111111111101;
			7'b1010000: Y = 33'b000001111111111111111111111111110;
			7'b1010001: Y = 33'b000001111111111111111111111111111;
			7'b1010010: Y = 33'b000011111111111111111111111111100;
			7'b1010011: Y = 33'b000011111111111111111111111111101;
			7'b1010100: Y = 33'b000011111111111111111111111111101;
			7'b1010101: Y = 33'b000011111111111111111111111111110;
			7'b1010110: Y = 33'b000011111111111111111111111111111;
			7'b1010111: Y = 33'b000111111111111111111111111111100;
			7'b1011000: Y = 33'b000111111111111111111111111111100;
			7'b1011001: Y = 33'b000111111111111111111111111111101;
			7'b1011010: Y = 33'b000111111111111111111111111111110;
			7'b1011011: Y = 33'b000111111111111111111111111111110;
			7'b1011100: Y = 33'b000111111111111111111111111111111;
			7'b1011101: Y = 33'b001111111111111111111111111111100;
			7'b1011110: Y = 33'b001111111111111111111111111111100;
			7'b1011111: Y = 33'b001111111111111111111111111111101;
			7'b1100000: Y = 33'b001111111111111111111111111111110;
			7'b1100001: Y = 33'b001111111111111111111111111111110;
			7'b1100010: Y = 33'b001111111111111111111111111111111;
			7'b1100011: Y = 33'b001111111111111111111111111111111;
			7'b1100100: Y = 33'b011111111111111111111111111111100;
			7'b1100101: Y = 33'b011111111111111111111111111111100;
			7'b1100110: Y = 33'b011111111111111111111111111111101;
			7'b1100111: Y = 33'b011111111111111111111111111111101;
			7'b1101000: Y = 33'b011111111111111111111111111111110;
			7'b1101001: Y = 33'b011111111111111111111111111111110;
			7'b1101010: Y = 33'b011111111111111111111111111111111;
			7'b1101011: Y = 33'b011111111111111111111111111111111;
			7'b1101100: Y = 33'b011111111111111111111111111111111;
			7'b1101101: Y = 33'b111111111111111111111111111111100;
			7'b1101110: Y = 33'b111111111111111111111111111111100;
			7'b1101111: Y = 33'b111111111111111111111111111111100;
			7'b1110000: Y = 33'b111111111111111111111111111111101;
			7'b1110001: Y = 33'b111111111111111111111111111111101;
			7'b1110010: Y = 33'b111111111111111111111111111111101;
			7'b1110011: Y = 33'b111111111111111111111111111111110;
			7'b1110100: Y = 33'b111111111111111111111111111111110;
			7'b1110101: Y = 33'b111111111111111111111111111111110;
			7'b1110110: Y = 33'b111111111111111111111111111111110;
			7'b1110111: Y = 33'b111111111111111111111111111111110;
			7'b1111000: Y = 33'b111111111111111111111111111111110;
			7'b1111001: Y = 33'b111111111111111111111111111111111;
			7'b1111010: Y = 33'b111111111111111111111111111111111;
			7'b1111011: Y = 33'b111111111111111111111111111111111;
			7'b1111100: Y = 33'b111111111111111111111111111111111;
			7'b1111101: Y = 33'b111111111111111111111111111111111;
			7'b1111110: Y = 33'b111111111111111111111111111111111;
			7'b1111111: Y = 33'b111111111111111111111111111111111;
//			default: Y = 33'b000000000000000000000000000000000;
		endcase
	end
endmodule

